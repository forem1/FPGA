module top
(
    input             clk, rst, btn1, btn2, btn3, btn4, led1, led2, led3, led4
);

    always @ (posedge clk or posedge rst)
    begin
        //if (rst)
        //begin
        //end
        
    end

endmodule
